netcdf struct_3d_json_export_null_nodata {
dimensions:
	time = 3 ;
	lat = 10 ;
	lon = 5 ;
variables:
	short tos1(time, lat, lon) ;
		tos1:valid_min = -32768s ;
		tos1:valid_max = 32767s ;
		tos1:missing_value = 120s ;
		tos1:_FillValue = 120s ;
		tos1:cell_methods = "time: mean (interval: 30 minutes)" ;
		tos1:history = " At 16:37:23 on 01/11/2005: CMOR altered the data in the following ways: added 2.73150E+02 to yield output units; Cyclical dimension was output starting at a different lon;" ;
		tos1:long_name = "Sea Surface Temperature" ;
		tos1:original_name = "sosstsst" ;
		tos1:original_units = "degC" ;
		tos1:standard_name = "sea_surface_temperature" ;
		tos1:units = "K" ;
	short tos2(time, lat, lon) ;
		tos2:valid_min = -32768s ;
		tos2:valid_max = 32767s ;
		tos2:missing_value = 200s ;
		tos2:_FillValue = 200s ;
		tos2:cell_methods = "time: mean (interval: 30 minutes)" ;
		tos2:history = " At 16:37:23 on 01/11/2005: CMOR altered the data in the following ways: added 2.73150E+02 to yield output units; Cyclical dimension was output starting at a different lon;" ;
		tos2:long_name = "Sea Surface Temperature" ;
		tos2:original_name = "sosstsst" ;
		tos2:original_units = "degC" ;
		tos2:standard_name = "sea_surface_temperature" ;
		tos2:units = "K" ;
	double lat(lat) ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
		lat:long_name = "latitude" ;
		lat:original_units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
	double lon(lon) ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
		lon:long_name = "longitude" ;
		lon:original_units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:calendar = "360_day" ;
		time:long_name = "time" ;
		time:original_units = "seconds since 2001-1-1" ;
		time:standard_name = "time" ;
		time:units = "days since 2001-1-1" ;

// global attributes:
		:Conventions = "CF-1.0" ;
		:cmor_version = 0.96 ;
		:comment = "Test drive" ;
		:contact = "Sebastien Denvil, sebastien.denvil@ipsl.jussieu.fr" ;
		:experiment_id = "SRES A2 experiment" ;
		:history = "YYYY/MM/JJ: data generated; YYYY/MM/JJ+1 data transformed At 16:37:23 on 01/11/2005, CMOR rewrote data to comply with CF standards and IPCC Fourth Assessment requirements" ;
		:institution = "IPSL (Institut Pierre Simon Laplace, Paris, France)" ;
		:project_id = "IPCC Fourth Assessment" ;
		:realization = 1L ;
		:references = "Dufresne et al, Journal of Climate, 2015, vol XX, p 136" ;
		:source = "IPSL-CM4_v1 (2003) : atmosphere : LMDZ (IPSL-CM4_IPCC, 96x71x19), ocean ORCA2 (ipsl_cm4_v1_8, 2x2L31); sea ice LIM (ipsl_cm4_v" ;
		:table_id = "Table O1 (13 November 2004)" ;
		:title = "IPSL model output prepared for IPCC Fourth Assessment SRES A2 experiment" ;
data:

 tos1 =
  1, 2, 3, 4, 5,
  6, 7, 8, 9, 10,
  11, 12, 13, 14, 15,
  16, 17, 18, 19, 20,
  21, 22, 23, 24, 25,
  26, 27, 28, 29, 30,
  31, 32, 33, 34, 35,
  36, 37, 38, 39, 40,
  41, 42, 43, 44, 45,
  46, 47, 48, 49, 50,
  51, 52, 53, 54, 55,
  56, 57, 58, 59, 60,
  61, 62, 63, 64, 65,
  66, 67, 68, 69, 70,
  71, 72, 73, 74, 75,
  76, 77, 78, 79, 80,
  81, 82, 83, 84, 85,
  86, 87, 88, 89, 90,
  91, 92, 93, 94, 95,
  96, 97, 98, 99, 100,
  101, 102, 103, 104, 105,
  106, 107, 108, 109, 110,
  111, 112, 113, 114, 115,
  116, 117, 118, 119, _,
  121, 122, 123, 124, 125,
  126, 127, 128, 129, 130,
  131, 132, 133, 134, 135,
  136, 137, 138, 139, 140,
  141, 142, 143, 144, 145,
  146, 147, 148, 149, 150 ;

 tos2 =
  151, 152, 153, 154, 155,
  156, 157, 158, 159, 160,
  161, 162, 163, 164, 165,
  166, 167, 168, 169, 170,
  171, 172, 173, 174, 175,
  176, 177, 178, 179, 180,
  181, 182, 183, 184, 185,
  186, 187, 188, 189, 190,
  191, 192, 193, 194, 195,
  196, 197, 198, 199, _,
  201, 202, 203, 204, 205,
  206, 207, 208, 209, 210,
  211, 212, 213, 214, 215,
  216, 217, 218, 219, 220,
  221, 222, 223, 224, 225,
  226, 227, 228, 229, 230,
  231, 232, 233, 234, 235,
  236, 237, 238, 239, 240,
  241, 242, 243, 244, 245,
  246, 247, 248, 249, 250,
  251, 252, 253, 254, 255,
  256, 257, 258, 259, 260,
  261, 262, 263, 264, 265,
  266, 267, 268, 269, 270,
  271, 272, 273, 274, 275,
  276, 277, 278, 279, 280,
  281, 282, 283, 284, 285,
  286, 287, 288, 289, 290,
  291, 292, 293, 294, 295,
  296, 297, 298, 299, 300 ;

 lat = -79.5, -78.5, -77.5, -76.5, -75.5, -74.5, -73.5, -72.5, -71.5, -70.5 ;

 lon = 1, 3, 5, 7, 9 ;

 time = 15, 45, 0 ;
}
